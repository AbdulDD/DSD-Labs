`timescale 1ns / 1ps                // Compilation/simulation directive

module OnetoFourDemultiplexer(input S1, S0, D, output Y[3:0]);

// Assign statement
assign 


endmodule
